module full_addr(

);

endmodule 