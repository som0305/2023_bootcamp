module testbench();

reg [31:0] a;
reg [31:0] b;
reg cin;
wire [31:0] sum;
wire cout;


