module CLA_32bit(
    input [31:0] a, b,
    input cin,
    output [31:0] sum,
    output cout
);

wire [2:0] carry;







