module testbench();
