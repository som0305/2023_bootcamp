module CL_32bit(
    input [31:0] a, b,
    input cin,
    output [31:0] sum,
    output cout
);

wire carry;

